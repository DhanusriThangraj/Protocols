VCD info: dumpfile Waves.vcd opened for output.
VCD warning: $dumpvars: Package ($unit) is not dumpable with VCD.
---WRITE--- Addr=a Data=aaaa
---WRITE--- Addr=b Data=bbbb
---WRITE--- Addr=c Data=cccc
---READ---  Addr=a Data=aaaa
---READ---  Addr=b Data=bbbb
---READ---  Addr=c Data=cccc
testbench.sv:51: $finish called at 355 (1s)
Finding VCD file...
./Waves.vcd
[2025-08-22 13:00:07 UTC] Opening EPWave...
Done
